module sam_nand2(a,b,c);
input a,b;
output c;
nand n2(c,a,b);
endmodule 

